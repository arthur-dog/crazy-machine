library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.utils.all;

entity section_2_b is
    port (
        clk_in : in std_logic;
        reset : in std_logic;


    )
end section_2_b;

architecture base of section_2_b is
begin
end base;
