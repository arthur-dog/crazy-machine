library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity servo_test_leds is
    Port (
        clk_50MHz : in  STD_LOGIC;      -- 50 MHz clock
        sw0       : in  STD_LOGIC;      -- Position select (mid = 45°)
        sw1       : in  STD_LOGIC;      -- Position select (max = 90°)
        led0      : out STD_LOGIC;      -- LED for SW0 (LEDR0)
        led1      : out STD_LOGIC;      -- LED for SW1 (LEDR1)
        servo_pwm : out STD_LOGIC       -- PWM output to servo
    );
end servo_test_leds;

architecture Behavioral of servo_test_leds is

    -- PWM timing constants
    constant PWM_PERIOD      : integer := 1000000;  -- 20ms = 1,000,000 @ 50MHz
    constant PULSE_0_DEG     : integer := 50000;    -- 1ms pulse = 0°
    constant PULSE_45_DEG    : integer := 75000;    -- 1.25ms pulse = ~45°
    constant PULSE_90_DEG    : integer := 100000;    -- 1.5ms pulse = ~90°

    signal counter      : integer range 0 to PWM_PERIOD := 0;
    signal pulse_width  : integer := PULSE_0_DEG;
    signal pwm_out      : std_logic := '0';

begin

    -- PWM signal generation
    process(clk_50MHz)
    begin
        if rising_edge(clk_50MHz) then
            -- Determine pulse width based on switches
            if sw1 = '1' then
                pulse_width <= PULSE_90_DEG;  -- Max = 90°
            elsif sw0 = '1' then
                pulse_width <= PULSE_45_DEG;  -- Mid = ~45°
            else
                pulse_width <= PULSE_0_DEG;   -- Min = 0°
            end if;

            -- PWM counter
            if counter < PWM_PERIOD then
                counter <= counter + 1;
            else
                counter <= 0;
            end if;

            -- PWM signal output
            if counter < pulse_width then
                pwm_out <= '1';
            else
                pwm_out <= '0';
            end if;
        end if;
    end process;

    -- Assign LEDs to match switch state
    led0 <= sw0;
    led1 <= sw1;

    -- Assign final PWM output
    servo_pwm <= pwm_out;

end Behavioral;
